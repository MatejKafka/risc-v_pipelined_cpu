`ifndef PACKAGE_TYPES
`define PACKAGE_TYPES

typedef logic [31:0] Reg;
`define REG_ADDRESS_WIDTH 5
typedef logic [`REG_ADDRESS_WIDTH-1:0] RegAddress;

`endif